`include "Opcode.vh"

module mmio (
    input clk,
    input [31:0] instr,
    input [31:0] pc_wb,
    input [31:0] instr_ex,
    input [31:0] instr_wb,
    input [31:0] alu_out,
    input [31:0] alu_reg_out
);



endmodule