`include "Opcode.vh"

module branch_predictor (
    output branch_taken
);
    
    assign branch_taken = 1;
endmodule